class mx_sequencer extends uvm_sequencer#(seqitem);
  `uvm_component_utils(mx_sequencer)
  
  
  function new(string name="mx_sequencer", uvm_component parent);
    super.new(name,parent);
  endfunction
  
  
  
  
  
endclass
